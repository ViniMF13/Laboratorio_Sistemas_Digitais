LIBRARY ieee;
USE ieee.std_logic_1164.all;

entity fulladder is
    port ( 
		  Cin : in std_logic;
		  x   : in std_logic;
		  y   : in std_logic;
		  s   : out std_logic;
		  Cout : out std_logic
        );
end fulladder;
architecture RTL OF fulladder is
begin
    s <= x XOR y XOR Cin;
    Cout <= (x AND y) OR (Cin AND x) OR (Cin AND y);
end RTL ;